*** SPICE deck for cell VCOSim{sch} from library VCO
*** Created on Tue Mar 18, 2025 10:29:18
*** Last revised on Tue Mar 18, 2025 12:44:11
*** Written on Tue Mar 18, 2025 12:44:19 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT VCO__NOT FROM CELL NOT{sch}
.SUBCKT VCO__NOT A Y
** GLOBAL gnd
** GLOBAL vdd
MM1 Y A vdd vdd PMOS L=0.2U W=2U
MM2 Y A gnd gnd NMOS L=0.2U W=1U
.ENDS VCO__NOT

.global gnd vdd

*** TOP LEVEL CELL: VCOSim{sch}
XN1 Y net@1 VCO__NOT
XN2 net@1 net@2 VCO__NOT
XN3 net@2 Y VCO__NOT

* Spice Code nodes in cell cell 'VCOSim{sch}'
.include ../180nm.lib
vdd vdd 0 1.8
.ic v(Y)=.1
.control
tran 0.1p 1000p
plot v(Y)
.endc
.end
.END
